// this is test file
module moduleName (
    ports
);
    
endmodule